// Предсказатель переходов

// Позволяет ускорить работу программы при выполнении циклов
// и операторов ветвления, в которых проверяемое условие чаще
// истинное, чем ложное

module branch_predictor
(
	input  wire [31:0] instr,
	input  wire [31:0] instr_addr,

	output wire [31:0] next_addr
);

wire [31:0] j_imm = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
wire [31:0] b_imm = {{20{instr[31]}}, instr[7], instr[30:25], instr[11:8], 1'b0};

assign next_addr =

        // Если это JAL, то сразу выбрать инструкцию по адресу перехода
	instr[6:0] == 7'h6F ? instr_addr + j_imm :

	// Если это Bxx и переход выполняется назад, то выбрать инструкцию
	// по адресу перехода, чтобы цикл выполнялся быстрее (случай do ... while)
	// Если это Bxx и переход выполняется вперёд, то выбрать следующую
	// инструкцию, чтобы оператор if выполнялся быстрее (случай if ... else)
	instr[6:0] == 7'h63 && instr[31] ? instr_addr + b_imm :

	// Если ни одно условие не сработало, то выбрать следующую инструкцию
	instr_addr + 3'd4;

endmodule
